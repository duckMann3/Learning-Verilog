module hello;
  initial
    begin
      $display("Hello Wolrd!");
      $finish;
    end
endmodule
